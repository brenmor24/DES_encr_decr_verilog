module encrypt_value(
input [63:0]key,
input [63:0]value,
output reg [63:0]msg
);

endmodule
